CIRCUIT Example.msk
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
Vb 7 0 PULSE(0.00 1.20 0.48N 0.03N 0.03N 0.48N 1.00N)
Va 8 0 PULSE(0.00 1.20 0.23N 0.03N 0.03N 0.23N 0.50N)
*
* List of nodes
* "and" corresponds to n�3
* "N5" corresponds to n�5
* "N6" corresponds to n�6
* "b" corresponds to n�7
* "a" corresponds to n�8
* "N9" corresponds to n�9
*
* MOS devices
MN1 0 5 3 0 N1  W= 0.24U L= 0.12U
MN2 6 7 5 0 N1  W= 0.24U L= 0.12U
MN3 0 8 6 0 N1  W= 0.24U L= 0.12U
MP1 1 5 3 1 P1  W= 0.72U L= 0.12U
MP2 5 7 1 1 P1  W= 0.72U L= 0.12U
MP3 1 8 5 1 P1  W= 0.72U L= 0.12U
*
C2 1 0  2.615fF
C3 3 0  0.694fF
C5 5 0  0.706fF
C6 6 0  0.090fF
C7 7 0  0.314fF
C8 8 0  0.314fF
C9 9 0  0.443fF
*
* Extra RLC
*
Radd1 3 9 5
*
*
* n-MOS BSIM4 :
* low leakage
.MODEL N1 NMOS LEVEL=14 VTO=0.40 U0=0.050 TOX= 2.0E-9 LINT=0.010U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.540 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.6 U0=0.050 UA=3.000e-15
+WINT=0.020U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.050
+XJ=0.150U NDEP=170.000e15 PCLM=1.100
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS BSIM4:
* low leakage
.MODEL P1 PMOS LEVEL=14 VTO=-0.45 U0=0.018 TOX= 2.0E-9 LINT=0.010U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.540 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.6 U0=0.018 UA=1.500e-15
+WINT=0.020U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.050
+XJ=0.150U NDEP=170.000e15 PCLM=0.700
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.TRAN 0.1N 2.00N
* (Pspice)
.PROBE
.END
