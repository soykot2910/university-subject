CIRCUIT C:\Users\Sk Buland\Downloads\MICROWIND_3.1\examples\Nand2.MSK
*
* IC Technology: CMOS 90nm, 6 Metal Copper - strained SiGe - LowK
*
VDD 1 0 DC 1.20
Va 6 0 DC 0 PULSE(0.00 1.20 0.23N 0.02N 0.02N 0.23N 0.50N)
Vb 7 0 DC 0 PULSE(0.00 1.20 0.48N 0.02N 0.02N 0.48N 1.00N)
*
* List of nodes
* "nand2" corresponds to n�3
* "N5" corresponds to n�5
* "a" corresponds to n�6
* "b" corresponds to n�7
*
* MOS devices
MN1 5 7 3 0 N1  W= 0.20U L= 0.10U
MN2 0 6 5 0 N1  W= 0.20U L= 0.10U
MP1 3 7 1 1 P1  W= 0.60U L= 0.10U
MP2 1 6 3 1 P1  W= 0.60U L= 0.10U
*
C2 1 0  1.518fF
C3 3 0  0.658fF
C5 5 0  0.071fF
C6 6 0  0.149fF
C7 7 0  0.149fF
*
*
* n-MOS BSIM4 :
* low leakage
.MODEL N1 NMOS LEVEL=14 VTHO=0.28 U0=0.060 TOXE= 1.2E-9 LINT=0.015U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.570 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  0.9 U0=0.060 UA=3.400e-15
+WINT=0.005U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.010
+XJ=0.150U NDEP=170.000e15 PCLM=1.100
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* p-MOS BSIM4:
* low leakage
.MODEL P1 PMOS LEVEL=14 VTHO=-0.32 U0=0.027 TOXE= 1.2E-9 LINT=0.015U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.570 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.9 U0=0.027 UA=2.200e-15
+WINT=0.005U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.010
+XJ=0.150U NDEP=170.000e15 PCLM=0.700
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* Transient analysis
*
* (Winspice)
.options temp=27.0
.control
tran 0.1N 2.00N
print  V(6) V(3) V(7) > out.txt
plot  V(6) V(3) V(7)
.endc
.END
